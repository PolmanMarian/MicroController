library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Program_rom is
	port(
	adress : in std_logic_vector(7 downto 0) := "00000000"; --adresa default cand incepe programul este 0
	instruction : out std_logic_vector(15 downto 0) := "1111111111111111"; --codificarea instructiunii care nu face nimic
	clock : in std_logic;
	enable : in std_logic
	);
end Program_rom;

architecture Behavioral of Program_rom is
type rom_array is array (0 to 255) of std_logic_vector(15 downto 0);
constant rom : rom_array :=(
"0100000111111010",--00 ADD S1,FAx;
"0000010110011000",--01 Load S5,98x;
"0000110000011010",--02 Load SC,1Ax;
"1100000111000001",--03 And S1,SC;
"1100001011110000",--04 Load S2,SF;
"0100000111000000",--05 ADD S1,C0x;
"1001110000000101",--06 JMPNC 05x;
"1100110001010101",--07 ADDCY SC,S5;
"0011011011100011",--08 XOR S6,E3;
"1100001101010010",--09 OR S3,S5;
"0110010001000100",--0A SUB S4,44x;
"1100011001000111",--0B SUBCY S6,S4;
"1100100010010100",--0C ADD S8,S9;
"1001000000001111",--0D JUMPZ 0F;
"0010011111110101",--0E OR S7,F5;
"0101100111101110",--0F ADD S9,EE;
"1001110000001100",--10 JUMPNC 0Cx;
"1111111111111111",--HOOO
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
"0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000");
begin
	process(clock , adress , enable)
	begin
		if enable = '1' then
			if rising_edge(clock) then
				instruction <= rom(to_integer(unsigned(adress)));
			end if;
		end if;
	end process;
end architecture;

